library verilog;
use verilog.vl_types.all;
entity g06_lab2_vlg_vec_tst is
end g06_lab2_vlg_vec_tst;
