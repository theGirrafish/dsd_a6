library verilog;
use verilog.vl_types.all;
entity gA6_lab3_vlg_vec_tst is
end gA6_lab3_vlg_vec_tst;
