library verilog;
use verilog.vl_types.all;
entity gA6_block_blackjack_vlg_vec_tst is
end gA6_block_blackjack_vlg_vec_tst;
