library verilog;
use verilog.vl_types.all;
entity Block2_vlg_vec_tst is
end Block2_vlg_vec_tst;
