library verilog;
use verilog.vl_types.all;
entity gA6_lab4_vlg_check_tst is
    port(
        ace_out         : in     vl_logic;
        legal_play      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gA6_lab4_vlg_check_tst;
